module main

struct OpenApi {
	
}