module open_api

import x.json2 { Any }
import json

struct RequestBody {
pub mut:
	description string
	content     map[string]MediaType
	required    bool
}

pub fn (mut request_body RequestBody) from_json(json Any) ? {
	object := json.as_map()
	check_required<RequestBody>(object, 'content') ?

	for key, value in object {
		match key {
			'description' {
				request_body.description = value.str()
			}
			'content' {
				request_body.content = decode_map<MediaType>(value.json_str()) or {
					return error('Failed RequestBody decoding: $err')
				}
			}
			'required' {
				request_body.required = value.bool()
			}
			else {}
		}
	}
}
